library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity DO5 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_DO5 of DO5 is
begin
	y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000001111110000000001000000100000001000000010000011111111111111111111111111111111001000000010000000010000010000000000111110000000000000000000000000000000000000000000000000000000";

end architecture; 










--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000111111000000
--0001000000100000
--0010000000100000
--1111111111111111
--1111111111111111
--0010000000100000
--0001000001000000
--0000111110000000
--0000000000000000
--0000000000000000
--0000000000000000



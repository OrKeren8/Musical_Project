library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity si1_1 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_si1_1 of si1_1 is
begin
	
y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111110000000001111111100000111111111111111111111111111111110001111111100000000111111100000000011111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";


	end architecture;

--y<="0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000011110000000
--0000111111000000
--0001111111100000
--1111111111111111
--1111111111111111
--0001111111100000
--0001111111000000
--0001111110000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000";

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity SOL1 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_SOL1 of SOL1 is
begin
	y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000011111100000000011111110000000011111111000011111111111111111111111111111111000011111111000000000111111000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		

end architecture; 





--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000001111110000
--0000011111110000
--0000111111110000
--1111111111111111
--1111111111111111
--0000111111110000
--0000011111100000
--0000001111000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000






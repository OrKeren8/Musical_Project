library ieee;
use ieee.std_logic_1164.all;

package Notes is

constant do1 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000111111100000000111111110000000111111111000001111111111111000111111111111100000111111111000000011111111100000000111111100000000001111100000000000000000000000000000000000000";


--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000011111110000
--0000111111110000
--0001111111110000
--0111111111111100
--0111111111111100
--0001111111110000
--0000111111100000
--0000011111000000
--0000000000000000
--0000000000000000
--0000000000000000

constant do2 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000111111100000000110000011000000110000001100001111111111111000111111111111100000110000001100000011000000110000000110000110000000001111100000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000011111110000
--0000110000011000
--0001100000011000
--0111111111111100
--0111111111111100
--0001100000011000
--0001100000011000
--0000110000110000
--0000011111000000
--0000000000000000
--0000000000000000

constant do3 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000001100000000000000110000000000000011110000000000001111000000000000111111000000000011111100000000001100111000000000110011111111111111111111111111111111111000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000000011000000000000001100000000000000110000000001111111000000001111111100000001111111110000011111111111110001111111111111000001111111110000000111111111000000001111111000000000011111000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001111000
--0000000001111000
--0000000001111110
--0000000001111110
--0000000001100111
--0000000001100111
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001100000
--0000111111100000
--0001111111100000
--0011111111100000
--1111111111111000
--1111111111111000
--0011111111100000
--0011111111100000
--0001111111000000
--0000111110000000
--0000000000000000
--0000000000000000

constant do4 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000001100000000000000110000000000000011110000000000001111000000000000111111000000000011111100000000001100111000000000110011111111111111111111111111111111111000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000000011000000000000001100000000000000110000000001111111000000001111111100000001111111110000011111111111110001111111111111000001111111110000000111111111000000001111111000000000011111000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001111000
--0000000001111000
--0000000001111110
--0000000001111110
--0000000001100111
--0000000001100111
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001100000
--0000111111100000
--0001111111100000
--0011111111100000
--1111111111111000
--1111111111111000
--0011111111100000
--0011111111100000
--0001111111000000
--0000111110000000
--0000000000000000
--0000000000000000

constant do5 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000001111110000000001000000100000001000000010000011111111111111111111111111111111001000000010000000010000010000000000111110000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000111111000000
--0001000000100000
--0010000000100000
--1111111111111111
--1111111111111111
--0010000000100000
--0001000001000000
--0000111110000000
--0000000000000000
--0000000000000000
--0000000000000000

constant re1 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000111111111111111111111111111111110000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000111111000000000111111100000000111111110000000011111111000000001111111100000000111111110000000001111110000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
--	   0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		1111111111111111
--		1111111111111111
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		1111111111111111
--		1111111111111111
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		1111111111111111
--		1111111111111111
--		0000011111100000
--		0000111111100000
--		0001111111100000
--		0001111111100000
--		0001111111100000
--		0001111111100000
--		0000111111000000
--		0000011110000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000"; 

constant re2 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000111111111111111111111111111111110000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000111111000000000100001100000000100000110000000010000011000000001000001100000000100000110000000001000010000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 

--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		1111111111111111
--		1111111111111111
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		1111111111111111
--		1111111111111111
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		0000000001100000
--		1111111111111111
--		1111111111111111
--		0000011111100000
--		0000100001100000
--		0001000001100000
--		0001000001100000
--		0001000001100000
--		0001000001100000
--		0000100001000000
--		0000011110000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant re3 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000111100000000000011110000111111111111111111111111111111110000000011001110000000001100111000000000110000100000000011000010000000001100000000000000110000000000000011000000000000001100000011111111111111111111111111111111000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000001111111111111111111111111111111100011111110000000011111111000000001111111100000000111111110000000011111111000000000111111000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

constant re4 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000111100000000000011110000111111111111111111111111111111110000000011001110000000001100111000000000110000100000000011000010000000001111000000000000111100000000000011111100000000001111110011111111111111111111111111111111000000001100001000000000110000100000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000001111111111111111111111111111111100011111110000000011111111000000001111111100000000111111110000000011111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

constant re5 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100001111110000000001000001000000001000000100000000100000010000000010000001000000001000000100000000010000100000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--    0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000111111000000
--		0001000001000000
--		0010000001000000
--		0010000001000000
--		0010000001000000
--		0010000001000000
--		0001000010000000
--		0000111100000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant mi1 : std_logic_vector(0 to 1023) :=  "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000001111110000000001111111000000001111111100001111111111111111111111111111111100001111111100000000011111100000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000001111110000
--0000011111110000
--0000111111110000
--1111111111111111
--1111111111111111
--0000111111110000
--0000011111100000
--0000001111000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000


constant mi2 : std_logic_vector (0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000001111110000000001000011000000001000001100001111111111111111111111111111111100001000001100000000010000110000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000001111110000
--0000010000110000
--0000100000110000
--1111111111111111
--1111111111111111
--0000100000110000
--0000010000110000
--0000001111100000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant mi3 : std_logic_vector (0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000110000000000000011000000000000001111000000000000111100000000000011111100000000001111110000000000110011100000000011000110111111111111111111111111111111110000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000011111111111111111111111111111111000000001100000000000000110000000000000011000000000000001100000000000000110000000000111111000000000111111100000000111111110000001111111111111111111111111111111100111111110000000001111111000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011110000
--0000000011110000
--0000000011111100
--0000000011111100
--0000000011001110
--0000000011000110
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000111111000000
--0001111111000000
--0011111111000000
--1111111111111111
--1111111111111111
--0011111111000000
--0001111111000000
--0000111110000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant mi4 : std_logic_vector (0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000110000000000000011000000000000001111000000000000111100000000000011111100000000001111110000000000110011100000000011000110111111111111111111111111111111110000000011110000000000001111000000000000111111000000000011111100000000001100111000000000110011100000000011000010000000001100001011111111111111111111111111111111000000001100000000000000110000000000000011000000000000001100000000000000110000000000111111000000000111111100000000111111110000001111111111111111111111111111111100111111110000000001111111000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011110000
--0000000011110000
--0000000011111100
--0000000011111100
--0000000011001110
--0000000011000110
--1111111111111111
--1111111111111111
--0000000011110000
--0000000011110000
--0000000011111100
--0000000011111100
--0000000011001110
--0000000011001110
--0000000011000010
--0000000011000010
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000111111000000
--0001111111000000
--0011111111000000
--1111111111111111
--1111111111111111
--0011111111000000
--0001111111000000
--0000111110000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant mi5 : std_logic_vector (0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000001000010000000001000000100001111111111111111111111111111111100001000000100000000010000100000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000001111100000
--0000010000100000
--0000100000010000
--1111111111111111
--1111111111111111
--0000100000010000
--0000010000100000
--0000001111100000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant fa1 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000111111000000000111111100000000111111110000000011111111000000001111111100000000111111110000000001111110000000000011110000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000001111110000
--0000011111110000
--0000111111110000
--0000111111110000
--0000111111110000
--0000111111110000
--0000011111100000
--0000001111000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant fa2 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000111111000000000100001100000000100000110000000010000011000000001000001100000000100000110000000001000010000000000011110000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000001111110000
--0000010000110000
--0000100000110000
--0000100000110000
--0000100000110000
--0000100000110000
--0000010000100000
--0000001111000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant fa3 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000000011000000000000001100000000000000111100000000000011110000000000001111110000000000111111000000000011001110000000001100111111111111111111111111111111111110000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000001111110000000001111111000000001111111100000000111111110000000011111111000000001111111100000000011111100000000000111100000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001111000
--0000000001111000
--0000000001111110
--0000000001111110
--0000000001100111
--0000000001100111
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000011111100000
--0000111111100000
--0001111111100000
--0001111111100000
--0001111111100000
--0001111111100000
--0000111111000000
--0000011110000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant fa4 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011110001111111111111111111111111111111100000000011111100000000001100111000000000110011100000000011000010000000001100001000000000111100000000000011110000000000001111110111111111111111111111111111111110000000001100111000000000110000100000000011000010000000001100000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000001111110000000001111111000000001111111100000000111111110000000011111111000000001111111100000000011111100000000000111100000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000001100000
--0000000001100000
--0000000001111000
--1111111111111111
--1111111111111111
--0000000001111110
--0000000001100111
--0000000001100111
--0000000001100001
--0000000001100001
--0000000001111000
--0000000001111000
--0000000001111110
--1111111111111111
--1111111111111111
--0000000001100111
--0000000001100001
--0000000001100001
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000011111100000
--0000111111100000
--0001111111100000
--0001111111100000
--0001111111100000
--0001111111100000
--0000111111000000
--0000011110000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant fa5 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000111100000000000100001000000000100000010000000010000001000000001000000100000000100000010000000001000010000000000011110000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000001111000000
--0000010000100000
--0000100000010000
--0000100000010000
--0000100000010000
--0000100000010000
--0000010000100000
--0000001111000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
constant sol1 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000011111100000000011111110000000011111111000011111111111111111111111111111111000011111111000000000111111000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000001111110000
--0000011111110000
--0000111111110000
--1111111111111111
--1111111111111111
--0000111111110000
--0000011111100000
--0000001111000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant sol2 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000011111100000000010000110000000010000011000011111111111111111111111111111111000010000011000000000100001100000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000001111110000
--0000010000110000
--0000100000110000
--1111111111111111
--1111111111111111
--0000100000110000
--0000010000110000
--0000001111100000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant sol3 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000001100000000000000110000000000000011110000000000001111000000000000111111000000000011111100000000001100111000000000110001101111111111111111111111111111111100000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000111111111111111111111111111111110000000011000000000000001100000000000000110000000000000011000000000000001100000000001111110000000001111111000000001111111100000011111111111111111111111111111111001111111100000000011111110000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011110000
--0000000011110000
--0000000011111100
--0000000011111100
--0000000011001110
--0000000011000110
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000111111000000
--0001111111000000
--0011111111000000
--1111111111111111
--1111111111111111
--0011111111000000
--0001111111000000
--0000111110000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant sol4 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000001100000000000000110000000000000011110000000000001111000000000000111111000000000011111100000000001100111000000000110001101111111111111111111111111111111100000000111100000000000011110000000000001111110000000000111111000000000011001110000000001100111000000000110000100000000011000010111111111111111111111111111111110000000011000000000000001100000000000000110000000000000011000000000000001100000000001111110000000001111111000000001111111100000011111111111111111111111111111111001111111100000000011111110000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011110000
--0000000011110000
--0000000011111100
--0000000011111100
--0000000011001110
--0000000011000110
--1111111111111111
--1111111111111111
--0000000011110000
--0000000011110000
--0000000011111100
--0000000011111100
--0000000011001110
--0000000011001110
--0000000011000010
--0000000011000010
--1111111111111111
--1111111111111111
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000000011000000
--0000111111000000
--0001111111000000
--0011111111000000
--1111111111111111
--1111111111111111
--0011111111000000
--0001111111000000
--0000111110000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000 

constant sol5 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000010000100000000010000001000011111111111111111111111111111111000010000001000000000100001000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";		

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000001111100000
--0000010000100000
--0000100000010000
--1111111111111111
--1111111111111111
--0000100000010000
--0000010000100000
--0000001111100000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000

constant la1 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000111111111111111111111111111111110000011111100000000011111110000000011111111000000001111111100000000111111110000000011111111000000000111111000000000001111000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

	--	   0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		1111111111111111
	--		1111111111111111
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		1111111111111111
	--		1111111111111111
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		1111111111111111
	--		1111111111111111
	--		0000011111100000
	--		0000111111100000
	--		0001111111100000
	--		0001111111100000
	--		0001111111100000
	--		0001111111100000
	--		0000111111000000
	--		0000011110000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000";
constant la2 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000111111111111111111111111111111110000011111100000000010000110000000010000011000000001000001100000000100000110000000010000011000000000100001000000000001111000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--	y<="	0000000000000000
--			0000000000000000
--			0000000000000000
--			0000000000000000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		1111111111111111
	--		1111111111111111
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		1111111111111111
	--		1111111111111111
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		0000000001100000
	--		1111111111111111
	--		1111111111111111
	--		0000011111100000
	--		0000100001100000
	--		0001000001100000
	--		0001000001100000
	--		0001000001100000
	--		0001000001100000
	--		0000100001000000
	--		0000011110000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000";


constant la3 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011110000000000001111000011111111111111111111111111111111000000001100111000000000110011100000000011000010000000001100001000000000110000000000000011000000000000001100000000000000110000001111111111111111111111111111111100000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000111111111111111111111111111111110000111111000000000111111100000000111111110000000011111111000000001111111100000000111111110000000001111110000000000011110000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--	y<="	0000000000000000
--			0000000000000000
--			0000000000000000
--			0000000000000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011110000
	--		0000000011110000
	--		1111111111111111
	--		1111111111111111
	--		0000000011001110
	--		0000000011001110
	--		0000000011000010
	--		0000000011000010
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		1111111111111111
	--		1111111111111111
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		1111111111111111
	--		1111111111111111
	--		0000111111000000
	--		0001111111000000
	--		0011111111000000
	--		0011111111000000
	--		0011111111000000
	--		0011111111000000
	--		0001111110000000
	--		0000111100000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000";

constant la4 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011110000000000001111000011111111111111111111111111111111000000001100111000000000110011100000000011000010000000001100001000000000111100000000000011110000000000001111110000000000111111001111111111111111111111111111111100000000110000100000000011000010000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000111111111111111111111111111111110000111111000000000111111100000000111111110000000011111111000000001111111100000000111111110000000001111110000000000011110000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--	y<="	0000000000000000
--			0000000000000000
--			0000000000000000
--			0000000000000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011110000
	--		0000000011110000
	--		1111111111111111
	--		1111111111111111
	--		0000000011001110
	--		0000000011001110
	--		0000000011000010
	--		0000000011000010
	--		0000000011110000
	--		0000000011110000
	--		0000000011111100
	--		0000000011111100
	--		1111111111111111
	--		1111111111111111
	--		0000000011000010
	--		0000000011000010
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		1111111111111111
	--		1111111111111111
	--		0000111111000000
	--		0001111111000000
	--		0011111111000000
	--		0011111111000000
	--		0011111111000000
	--		0011111111000000
	--		0001111110000000
	--		0000111100000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000";

constant la5 : std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000111111000000000100000100000000100000010000000010000001000000001000000100000000100000010000000001000010000000000011110000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--	y<="	0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000111111000000
	--		0001000001000000
	--		0010000001000000
	--		0010000001000000
	--		0010000001000000
	--		0010000001000000
	--		0001000010000000
	--		0000111100000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000

	
constant si1 : std_logic_vector(0 to 1023) := "0000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000111111000000000111111100000000111111110000111111111111111111111111111111110000111111110000000001111110000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		1111111111111111
--		1111111111111111
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		1111111111111111
--		1111111111111111
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000001111110000
--		0000011111110000
--		0000111111110000
--		1111111111111111
--		1111111111111111
--		0000111111110000
--		0000011111100000
--		0000001111000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant si2 :std_logic_vector(0 to 1023) := "0000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000111111000000000100001100000000100000110000111111111111111111111111111111110000100000110000000001000110000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		1111111111111111
--		1111111111111111
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		1111111111111111
--		1111111111111111
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000000000110000
--		0000001111110000
--		0000010000110000
--		0000100000110000
--		1111111111111111
--		1111111111111111
--		0000100000110000
--		0000010001100000
--		0000001111000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant si3 :std_logic_vector(0 to 1023) := "0000000011000000000000001100000000000000111100000000000011110000000000001111110000000000111111000000000011001110000000001100111011111111111111111111111111111111000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000001111111111111111111111111111111100000000110000000000000011000000000000001100000000000000110000000000000011000000000011111100000000011111110000000011111111000000111111111111111111111111111111110011111111000000000111111000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--		0000000011000000
--		0000000011000000
--		0000000011110000
--		0000000011110000
--		0000000011111100
--		0000000011111100
--		0000000011001110
--		0000000011001110
--		1111111111111111
--		1111111111111111
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		1111111111111111
--		1111111111111111
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000111111000000
--		0001111111000000
--		0011111111000000
--		1111111111111111
--		1111111111111111
--		0011111111000000
--		0001111110000000
--		0000111100000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant si4 :std_logic_vector(0 to 1023) := "0000000011000000000000001100000000000000111100000000000011110000000000001111110000000000111111000000000011001110000000001100111011111111111111111111111111111111000000001111000000000000111100000000000011111100000000001111110000000000110011100000000011001110000000001100001000000000110000101111111111111111111111111111111100000000110000000000000011000000000000001100000000000000110000000000000011000000000011111100000000011111110000000011111111000000111111111111111111111111111111110011111111000000000111111000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--		0000000011000000
--		0000000011000000
--		0000000011110000
--		0000000011110000
--		0000000011111100
--		0000000011111100
--		0000000011001110
--		0000000011001110
--		1111111111111111
--		1111111111111111
--		0000000011110000
--		0000000011110000
--		0000000011111100
--		0000000011111100
--		0000000011001110
--		0000000011001110
--		0000000011000010
--		0000000011000010
--		1111111111111111
--		1111111111111111
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000000011000000
--		0000111111000000
--		0001111111000000
--		0011111111000000
--		1111111111111111
--		1111111111111111
--		0011111111000000
--		0001111110000000
--		0000111100000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant si5 :std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000010000010000000010000001000000111111111111111111111111111111110010000001000000000100001000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000111111000000
--		0001000001000000
--		0010000001000000
--		1111111111111111
--		1111111111111111
--		0010000001000000
--		0001000010000000
--		0000111100000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		1111111111111111
--		1111111111111111
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000
--		0000000000000000

constant do1_1 :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000111100000000000111111000000000111111110000000011111111000000001111111100000000111111110000000011111110000000001111110000000111111111111111111111111111111110001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--	y<="	0000000000000000
--			0000000000000000
--			0000000000000000
--			0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
--			0000000000000000
--			0000000000000000
--			0000000000000000
--			0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000011110000000
	--		0000111111000000
	--		0001111111100000
	--		0001111111100000
	--		0001111111100000
	--		0001111111100000
	--		0001111111000000
	--		0001111110000000
	--		1111111111111111
	--		1111111111111111
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		1111111111111111
	--		1111111111111111
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		1111111111111111
	--		1111111111111111
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0001100000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000";
--		


constant do1_2 :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000111100000000000100001000000000110000010000000011000001000000001100000100000000110000010000000011000010000000001111110000000111111111111111111111111111111110001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--y<="	0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000011110000000
--0000100001000000
--0001100000100000
--0001100000100000
--0001100000100000
--0001100000100000
--0001100001000000
--0001111110000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000";

constant do2_1 :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000111111100000000111111110000000111111111000001111111111111000111111111111100000111111111000000001111111000000000011111000000000000000000000000000000000000000000000000000000";


--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000111111
--1111111111111111
--1111111111111111
--0000000000111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000011111110000
--0000111111110000
--0001111111110000
--0111111111111100
--0111111111111100
--0001111111110000
--0000111111100000
--0000011111000000
--0000000000000000
--0000000000000000
--0000000000000000


constant do2_2 :std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000111111111111111111111111111111111111111111110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100001111111111111111111111111111111100000000001100000000000000110000000000000011000000000111111100000000111111110000000111111111000001111111111111000111111111111100000111111111000000001111111000000000011111000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111110000
--1111111111111111
--1111111111111111
--1111111111110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000011111110000
--0000111111110000
--0001111111110000
--0111111111111100
--0111111111111100
--0001111111110000
--0000111111100000
--0000011111000000
--0000000000000000
--0000000000000000
--0000000000000000

constant si2_1 :std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111110000000001111111100000111111111111111111111111111111110001111111100000000111111100000000011111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000000001111111111111000111111111111100011111111111110001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--y<="0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000011110000000
--0000111111000000
--0001111111100000
--1111111111111111
--1111111111111111
--0001111111100000
--0001111111000000
--0001111110000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001111111111111
--0001111111111111
--0001111111111111
--0001111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000";


constant si2_2 :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111110000000001111111100000111111111111111111111111111111110001111111100000000111111100000000011111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000001111100000000000111110000000000011111000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
--y<="0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000011110000000
--0000111111000000
--0001111111100000
--1111111111111111
--1111111111111111
--0001111111100000
--0001111111000000
--0001111110000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111100000000000
--1111100000000000
--1111100000000000
--1111100000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000";

constant si1_1 :std_logic_vector(0 to 1023) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111110000000001111111100000111111111111111111111111111111110001111111100000000111111100000000011111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--y<="0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000011110000000
--0000111111000000
--0001111111100000
--1111111111111111
--1111111111111111
--0001111111100000
--0001111111000000
--0001111110000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000";


constant si1_2 :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001000010000000001100000100000111111111111111111111111111111110001100000100000000110000100000000011111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000011111111111111111111111111111111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111111111111111111111111111111100011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--y<="0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000011110000000
--0000100001000000
--0001100000100000
--1111111111111111
--1111111111111111
--0001100000100000
--0001100001000000
--0001111110000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--1111111111111111
--1111111111111111
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0001100000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000";


constant lines :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000


constant shols :std_logic_vector(0 to 1023) :="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--y<="0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000


constant keySol :std_logic_vector(0 to 1023) :="0000000000111100000000001111111000000000100000010000000010000001000000011000000100000001100000010000000110000001000000011000000111111111111111111111111111111111000000011000000100000001100000010000000110000111000000011000011000000001100111000000000110011000000000011111000000000001111000001111111111111111111111111111111100000111100000000000011110000000000111011000000000011001100000000111000110000000011000011000000011000001100000001000000110000000111111111111111111111111111111111000000110000000100000011000000010000001100000001000000110000000100000011111100010000011111111001000011110000110100011011000001111111111111111111111111111111111110000011000001111000001100000110110000110000011001000011000001100110001100001100001000110001100000110011001100000001111111100001111111111111111111111111111111100000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000011001100000000011110110000000011111011000000001111101100000000111100110000000001100011000000000001001100000000000011110000000";

--Y=0000000000111100
--0000000011111110
--0000000010000001
--0000000010000001
--0000000110000001
--0000000110000001
--0000000110000001
--0000000110000001
--1111111111111111
--1111111111111111
--0000000110000001
--0000000110000001
--0000000110000111
--0000000110000110
--0000000110011100
--0000000110011000
--0000000111110000
--0000000111100000
--1111111111111111
--1111111111111111
--0000011110000000
--0000011110000000
--0001110110000000
--0001100110000000
--0111000110000000
--0110000110000000
--1100000110000000
--1000000110000000
--1111111111111111
--1111111111111111
--1000000110000000
--1000000110000000
--1000000110000000
--1000000110000000
--1000000111111000
--1000001111111100
--1000011110000110
--1000110110000011
--1111111111111111
--1111111111111111
--1100000110000011
--1100000110000011
--0110000110000011
--0010000110000011
--0011000110000110
--0001000110001100
--0001100110011000
--0000111111110000
--1111111111111111
--1111111111111111
--0000000110000000
--0000000110000000
--0000000110000000
--0000000110000000
--0000000110000000
--0000000110000000
--0001100110000000
--0011110110000000
--0111110110000000
--0111110110000000
--0111100110000000
--0011000110000000
--0000100110000000
--0000011110000000



type namesMatrix is array (127 downto 0) of std_logic_vector (1023 downto 0);
constant notesALL : namesMatrix :=
				(9=>do1, 10=>do2, 11=>do3, 12=>do4, 13=>do5, 
				17=>re1, 18=>re2, 19=>re3, 20=>re4, 21=>re5,
				25=>mi1, 26=>mi2, 27=>mi3, 28=>mi4, 29=>mi5,
				33=>fa1, 34=>fa2, 35=>fa3, 36=>fa4, 37=>fa5,
				41=>sol1, 42=>sol2, 43=>sol3, 44=>sol4, 45=>sol5,
				49=>la1, 50=>la2, 51=>la3, 52=>la4, 53=>la5,
				57=>si1, 58=>si2, 59=>si3, 60=>si4, 61=>si5,
				65=>do1_1, 66=>do1_2, 14=>do2_1,	15=>do2_2,
				105=>si1_1, 106=> si1_2, 110=>si2_1, 111=>si2_2,
				127=>lines, 0=>shols, 126=>keySol, 
				others=>shols														);


end package;



library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity PA3 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_PA3 of PA3 is
begin
	y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000001111111111111111111111111111111100000000011000000000000001100000000000000111100000000000011110000000000001111110000000000111111000000000011001110000000001100111111111111111111111111111111111110000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000011111111111111111111111111111111000001111110000000001111111000000001111111100000000111111110000000011111111000000001111111100000000011111100000000000111100000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
end architecture; 







--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001111000
--0000000001111000
--0000000001111110
--0000000001111110
--0000000001100111
--0000000001100111
--1111111111111111
--1111111111111111
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--0000000001100000
--1111111111111111
--1111111111111111
--0000011111100000
--0000111111100000
--0001111111100000
--0001111111100000
--0001111111100000
--0001111111100000
--0000111111000000
--0000011110000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000



library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity la4 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_la4 of la4 is
begin
	
y<="0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011110000000000001111000011111111111111111111111111111111000000001100111000000000110011100000000011000010000000001100001000000000111100000000000011110000000000001111110000000000111111001111111111111111111111111111111100000000110000100000000011000010000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000111111111111111111111111111111110000111111000000000111111100000000111111110000000011111111000000001111111100000000111111110000000001111110000000000011110000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

	end architecture;

--	y<="	0000000000000000
--			0000000000000000
--			0000000000000000
--			0000000000000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011110000
	--		0000000011110000
	--		1111111111111111
	--		1111111111111111
	--		0000000011001110
	--		0000000011001110
	--		0000000011000010
	--		0000000011000010
	--		0000000011110000
	--		0000000011110000
	--		0000000011111100
	--		0000000011111100
	--		1111111111111111
	--		1111111111111111
	--		0000000011000010
	--		0000000011000010
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		0000000011000000
	--		1111111111111111
	--		1111111111111111
	--		0000111111000000
	--		0001111111000000
	--		0011111111000000
	--		0011111111000000
	--		0011111111000000
	--		0011111111000000
	--		0001111110000000
	--		0000111100000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		1111111111111111
	--		1111111111111111
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000
	--		0000000000000000";
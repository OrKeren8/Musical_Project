library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package Melodies is

type matrix is array (255 downto 0) of std_logic_vector (6 downto 0);
constant keta0 : matrix := (

-------Little Yonatan----------

----------part 1---------------
	7 => "1111111",
	8  =>"1111110",  
	9  =>"1111111",  

	10  =>"0110001",  
	11  =>"0011001",  
	12  =>"0011010",  
	  13  =>"1111111",  

	  14  =>"0100001",  
	  15  =>"0010001",  
	  16  =>"0010010",  
	  17  =>"1111111",  

	  18  =>"0001001",  
	  19  =>"0010001",  
	  20  =>"0011001",  
	  21  =>"0100001",  
	  22  =>"0101001",  
	  23  =>"0101001",  
	  24  =>"0101010",  
	  25  =>"1111111",  

	  26  =>"0110001",  
	  27  =>"0011001",  
	  28  =>"0011010",  

	  29  =>"1111111",  
	  30  =>"1111111",  
	  31  =>"1111111",  
	  32  =>"1111111",  

-----part 2--------------
	  47  =>"1111111",  
	  48  =>"1111110",  
	  49  =>"1111111",  

	  50  =>"0100001",  
	  51  =>"0010001",  
	  52  =>"0010010",  
	  53  =>"1111111",  

	  54  =>"0001001",  
	  55  =>"0011001",  
	  56  =>"0101001",  
	  57  =>"0101001",  
	  58  =>"0001101",  
	  59  =>"1111111",  
	  60  =>"1111111",  
	  61  =>"1111111",  

	  62  =>"0010001",  
	  63  =>"0010001",  
	  64  =>"0010001",  
	  65  =>"0010001",  
	  66  =>"0010001",  
	  67  =>"0011001",  
	  68  =>"0100010",  

	  69  =>"1111111",  
	  70  =>"1111111",  
	  71  =>"1111111",  
	  72  =>"1111111",  

-----------part 3--------------

	  87  =>"1111111",  
	  88  =>"1111110",  
	  89  =>"1111111",  

	  90  =>"0011001",  
	  91  =>"0011001",  
	  92  =>"0011001",  
	  93  =>"0011001",  
	  94  =>"0011001",  
	  95  =>"0100001",  
	  96  =>"0101010",  
	  97  =>"1111111",  

	  98  =>"0110001",  
	  99  =>"0011001",  
	  100  =>"0011010",  
	  101  =>"1111111",  

	  102  =>"0100001",  
	  103  =>"0010001",  
	  104  =>"0010010",  
	  105  =>"1111111",  

	  106  =>"0001001",  
	  107  =>"0011001",  
	  108  =>"0101001",  
	  109  =>"0101001",  
	  110  =>"0001101",  

	  111  =>"1111111",  
	  112  =>"1111111",  

	 others => "0000000"
	);

constant keta1 : matrix := (
	 
-----"Uncle's Moshe farm"---

	
	9 =>"1111111",
	10 =>"1111110",
	11 =>"1111111",

	12 =>"0010001",
	13 =>"0101001",
	14 =>"0101001",
	15 =>"0101001",

	16 =>"0010001",
	17 =>"0011001",
	18 =>"0011001",
	19 =>"0010010",

	20 =>"1111111",
	21 =>"1101001",
	22 =>"1101001",
	23 =>"0110001",
	24 =>"0110001",
	25 =>"0101010",
	26 =>"1111111",
	27 =>"0010001",
	28 =>"1111111",
	29 =>"1111111",
	30 =>"1111111",

	 ---???2--

	49 =>"1111111",
	50 =>"1111110",
	51 =>"1111111",

	52 =>"1111111",
	53 =>"0101001",
	54 =>"0101001",
	55 =>"0101001",

	56 =>"0010001",
	57 =>"0011001",
	58 =>"0011001",
	59 =>"0010010",

	60 =>"1111111",
	61 =>"1101001",
	62 =>"1101001",
	63 =>"0110001",
	64 =>"0110001",
	65 =>"0101010",
	66 =>"1111111",
	67 =>"0010001",
	68 =>"1111111",
	69 =>"1111111",
	70 =>"1111111",

	----????--

	89 =>"1111111",
	90 =>"1111110",
	91 =>"1111111",

	92 =>"1111111",
	93 =>"0101001",
	94 =>"0101001",
	95 =>"0101001",
	96 =>"0010001",

	97 =>"0101001",
	98 =>"0101001",
	99 =>"0101010",

	100 =>"1111111",
	101 =>"0101001",
	102 =>"0101001",
	103 =>"0101001",
	104 =>"0010001",

	105 =>"0101001",
	106 =>"0101001",
	107 =>"0101001",
	108 =>"0010001",
	109 =>"1111111",
	110 =>"1111111",

	-----????--
	129 =>"1111111",
	130 =>"1111110",
	131 =>"1111111",

	132 =>"1111111",
	133 =>"0101001",
	134 =>"0101001",
	135 =>"0101001",

	136 =>"0010001",
	137 =>"0011001",
	138 =>"0011001",
	139 =>"0010010",

	140 =>"1111111",
	141 =>"1101001",
	142 =>"1101001",
	143 =>"0110001",
	144 =>"0110001",
	145 =>"0101101",
	146 =>"1111111",
	147 =>"1111111",
	148 =>"1111111",
	149 =>"1111111",
	150 =>"1111111",
	
	others => "0000000"
	);
	
constant keta2 : matrix := (


------Dear Mom----------
	
	
	0 => "0000000",
	10 => "1111111",
	11 => "1111110",
	12 => "1111111",
	
	13 => "0011001",
	14 => "0101001",
	15 => "0100001",
	16 => "0101001",
	
	17 => "0100010",
	18 => "1111111",

	19 => "0011010",
	20 => "1111111",
	
	21 => "0101010",
	22 => "1111111",
	
	23 => "0110010",
	24 => "1111111",
	
	25 => "0111101",
	26 => "1111111",
	27 => "1111111",
	28 => "1111111",
	29 => "1111111",

	 ---???2--
	50 => "1111111",
	51 => "1111110",
	52 => "1111111",
	
	53 => "1101001",
	54 => "1101001",
	55 => "1101001",
	
	56 => "0101001",
	57 => "0110001",
	58 => "0110001",

	59 => "0110010",
	60 => "1111111",
	
	61 => "0101001",
	62 => "0101001",
	63 => "0101001",
	64 => "0011001",
	
	65 => "0100001",
	66 => "0100001",
	67 => "0100001",
	68 => "0111001",
	69 => "1111111",

	----????--
	90 => "1111111",
	91 => "1111110",
	92 => "1111111",
	
	93 => "0101010",
	94 => "1111111",
	95 => "0100010",

	96 => "1111111",
	97 => "0011010",
	98 => "1111111",

	99 => "1101001",
	100 => "0101010",
	101 => "1111111",
	102 => "0100010",
	103 => "1111111",

	104 => "0011101",
	105 => "1111111",
	106 => "1111111",
	107 => "1111111",
	108 => "1111111",
	109 => "1111111",
	others => "0000000"
	);
--constant keta3 : matrix := ();
--constant keta4 : matrix := ();
--constant keta5 : matrix := ();
--constant keta6 : matrix := ();
--constant keta7 : matrix := ();

end package;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity keySol is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_keySol of keySol is
begin
		
	Y<="0000000000111100000000001111111000000000100000010000000010000001000000011000000100000001100000010000000110000001000000011000000111111111111111111111111111111111000000011000000100000001100000010000000110000111000000011000011000000001100111000000000110011000000000011111000000000001111000001111111111111111111111111111111100000111100000000000011110000000000111011000000000011001100000000111000110000000011000011000000011000001100000001000000110000000111111111111111111111111111111111000000110000000100000011000000010000001100000001000000110000000100000011111100010000011111111001000011110000110100011011000001111111111111111111111111111111111110000011000001111000001100000110110000110000011001000011000001100110001100001100001000110001100000110011001100000001111111100001111111111111111111111111111111100000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000011001100000000011110110000000011111011000000001111101100000000111100110000000001100011000000000001001100000000000011110000000";


end architecture; 








--Y=0000000000111100
--0000000011111110
--0000000010000001
--0000000010000001
--0000000110000001
--0000000110000001
--0000000110000001
--0000000110000001
--1111111111111111
--1111111111111111
--0000000110000001
--0000000110000001
--0000000110000111
--0000000110000110
--0000000110011100
--0000000110011000
--0000000111110000
--0000000111100000
--1111111111111111
--1111111111111111
--0000011110000000
--0000011110000000
--0001110110000000
--0001100110000000
--0111000110000000
--0110000110000000
--1100000110000000
--1000000110000000
--1111111111111111
--1111111111111111
--1000000110000000
--1000000110000000
--1000000110000000
--1000000110000000
--1000000111111000
--1000001111111100
--1000011110000110
--1000110110000011
--1111111111111111
--1111111111111111
--1100000110000011
--1100000110000011
--0110000110000011
--0010000110000011
--0011000110000110
--0001000110001100
--0001100110011000
--0000111111110000
--1111111111111111
--1111111111111111
--0000000110000000
--0000000110000000
--0000000110000000
--0000000110000000
--0000000110000000
--0000000110000000
--0001100110000000
--0011110110000000
--0111110110000000
--0111110110000000
--0111100110000000
--0011000110000000
--0000100110000000
--0000011110000000



library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package Melodies is

type matrix is array (255 downto 0) of std_logic_vector (6 downto 0);
constant keta0 : matrix := (

-------Little Yonatan----------
--keta0
----------part 1---------------
	7 => "1111111",
	8  =>"1111110",  
	9  =>"1111111",  

	10  =>"0110001",  
	11  =>"0011001",  
	12  =>"0011010",  
	13  =>"1111111",  

	14  =>"0100001",  
	15  =>"0010001",  
	16  =>"0010010",  
	17  =>"1111111",  

	18  =>"0001001",  
	19  =>"0010001",  
	20  =>"0011001",  
	21  =>"0100001",  
	22  =>"0101001",  
	23  =>"0101001",  
	24  =>"0101010",  
	25  =>"1111111",  

	26  =>"0110001",  
	27  =>"0011001",  
	28  =>"0011010",  

	29  =>"1111111",  
	30  =>"1111111",  
	31  =>"1111111",  
	32  =>"1111111",  

-----part 2--------------
	  47  =>"1111111",  
	  48  =>"1111110",  
	  49  =>"1111111",  

	  50  =>"0100001",  
	  51  =>"0010001",  
	  52  =>"0010010",  
	  53  =>"1111111",  

	  54  =>"0001001",  
	  55  =>"0011001",  
	  56  =>"0101001",  
	  57  =>"0101001",  
	  58  =>"0001101",  
	  59  =>"1111111",  
	  60  =>"1111111",  
	  61  =>"1111111",  

	  62  =>"0010001",  
	  63  =>"0010001",  
	  64  =>"0010001",  
	  65  =>"0010001",  
	  66  =>"0010001",  
	  67  =>"0011001",  
	  68  =>"0100010",  

	  69  =>"1111111",  
	  70  =>"1111111",  
	  71  =>"1111111",  
	  72  =>"1111111",  

-----------part 3--------------

	  87  =>"1111111",  
	  88  =>"1111110",  
	  89  =>"1111111",  

	  90  =>"0011001",  
	  91  =>"0011001",  
	  92  =>"0011001",  
	  93  =>"0011001",  
	  94  =>"0011001",  
	  95  =>"0100001",  
	  96  =>"0101010",  
	  97  =>"1111111",  

	  98  =>"0110001",  
	  99  =>"0011001",  
	  100  =>"0011010",  
	  101  =>"1111111",  

	  102  =>"0100001",  
	  103  =>"0010001",  
	  104  =>"0010010",  
	  105  =>"1111111",  

	  106  =>"0001001",  
	  107  =>"0011001",  
	  108  =>"0101001",  
	  109  =>"0101001",  
	  110  =>"0001101",  

	  111  =>"1111111",  
	  112  =>"1111111",  

	  others => "0000000"
	);

constant keta1 : matrix := (
	 
-----"Uncle's Moshe farm"---
--keta1
	
	9 =>"1111111",
	10 =>"1111110",
	11 =>"1111111",

	12 =>"0010001",
	13 =>"0101001",
	14 =>"0101001",
	15 =>"0101001",

	16 =>"0010001",
	17 =>"0011001",
	18 =>"0011001",
	19 =>"0010010",

	20 =>"1111111",
	21 =>"1101001",
	22 =>"1101001",
	23 =>"0110001",
	24 =>"0110001",
	25 =>"0101010",
	26 =>"1111111",
	27 =>"0010001",
	28 =>"1111111",
	29 =>"1111111",
	30 =>"1111111",

	 ---???2--

	49 =>"1111111",
	50 =>"1111110",
	51 =>"1111111",

	52 =>"1111111",
	53 =>"0101001",
	54 =>"0101001",
	55 =>"0101001",

	56 =>"0010001",
	57 =>"0011001",
	58 =>"0011001",
	59 =>"0010010",

	60 =>"1111111",
	61 =>"1101001",
	62 =>"1101001",
	63 =>"0110001",
	64 =>"0110001",
	65 =>"0101010",
	66 =>"1111111",
	67 =>"0010001",
	68 =>"1111111",
	69 =>"1111111",
	70 =>"1111111",

	----????--

	89 =>"1111111",
	90 =>"1111110",
	91 =>"1111111",

	92 =>"1111111",
	93 =>"0101001",
	94 =>"0101001",
	95 =>"0101001",
	96 =>"0010001",

	97 =>"0101001",
	98 =>"0101001",
	99 =>"0101010",

	100 =>"1111111",
	101 =>"0101001",
	102 =>"0101001",
	103 =>"0101001",
	104 =>"0010001",

	105 =>"0101001",
	106 =>"0101001",
	107 =>"0101001",
	108 =>"0010001",
	109 =>"1111111",
	110 =>"1111111",

	-----????--
	129 =>"1111111",
	130 =>"1111110",
	131 =>"1111111",

	132 =>"1111111",
	133 =>"0101001",
	134 =>"0101001",
	135 =>"0101001",

	136 =>"0010001",
	137 =>"0011001",
	138 =>"0011001",
	139 =>"0010010",

	140 =>"1111111",
	141 =>"1101001",
	142 =>"1101001",
	143 =>"0110001",
	144 =>"0110001",
	145 =>"0101101",
	146 =>"1111111",
	147 =>"1111111",
	148 =>"1111111",
	149 =>"1111111",
	150 =>"1111111",
	
	others => "0000000"
	);
	
constant keta2 : matrix := (


------Dear Mom----------
--keta2
--------part 1----------
	0 => "0000000",
	10 => "1111111",
	11 => "1111110",
	12 => "1111111",
	
	13 => "0011001",
	14 => "0101001",
	15 => "0100001",
	16 => "0101001",
	
	17 => "0100010",
	18 => "1111111",

	19 => "0011010",
	20 => "1111111",
	
	21 => "0101010",
	22 => "1111111",
	
	23 => "0110010",
	24 => "1111111",
	
	25 => "0111101",
	26 => "1111111",
	27 => "1111111",
	28 => "1111111",
	29 => "1111111",

--------part 2----------
	50 => "1111111",
	51 => "1111110",
	52 => "1111111",
	
	53 => "1101001",
	54 => "1101001",
	55 => "1101001",
	
	56 => "0101001",
	57 => "0110001",
	58 => "0110001",

	59 => "0110010",
	60 => "1111111",
	
	61 => "0101001",
	62 => "0101001",
	63 => "0101001",
	64 => "0011001",
	
	65 => "0100001",
	66 => "0100001",
	67 => "0100001",
	68 => "0111001",
	69 => "1111111",

--------part 3----------
	90 => "1111111",
	91 => "1111110",
	92 => "1111111",
	
	93 => "0101010",
	94 => "1111111",
	95 => "0100010",

	96 => "1111111",
	97 => "0011010",
	98 => "1111111",

	99 => "1101001",
	100 => "0101010",
	101 => "1111111",
	102 => "0100010",
	103 => "1111111",

	104 => "0011101",
	105 => "1111111",
	106 => "1111111",
	107 => "1111111",
	108 => "1111111",
	109 => "1111111",
	others => "0000000"
	);
	
constant keta3 : matrix := (
-------Happy Birthday----------
--keta3
----------part 1---------------
		10 => "1111111",
		11 => "1111110",
		12 => "1111111",
	
		13 => "0001110",
		14 => "0001111",
		15 => "0010001",
		16 => "0001001",	
		17 => "0100001",
	
		18 => "0011010",
		19 => "1111111",
		20 => "0001110",	
		21 => "0001111",
	
		22 => "0010001",	
		23 => "0001001",
		24 => "0101001",
	
		25 => "0100010",
		26 => "1111111",
		27 => "1111111",
		28 => "1111111",
		29 => "1111111",

----------part 2---------------

		50 => "1111111",
		51 => "1111110",
		52 => "1111111",
	
		53 => "0001110",
		54 => "0001111",
	
		55 => "1000001",	
		56 => "0110001",
		57 => "0100001",
	
		58 => "0011001",
		59 => "0010001",
		60 => "1101110",	
		61 => "1101111",
	
		62 => "0110001",
		63 => "0100001",
		64 => "0101001",
	
		65 => "0100010",
		66 => "1111111",
		67 => "1111111",
		68 => "1111111",
		69 => "1111111",
	others => "0000000"
	);
constant keta4 : matrix := (
-------Twinkle, Twinkle little star------------
--keta4
----------part 1---------------
		7 => "1111111",
		8 => "1111110",
		9 => "1111111",

		10 => "0001001",
		11 => "0001001",
		12 => "1111111",
		13 => "1111111",

		14 => "0101001",
		15 => "0101001",
		16 => "1111111",
		17 => "1111111",

		18 => "0110001",	
		19 => "1111111",
		20 => "0110001",
		21 => "1111111",
	
		22 => "1111111",
		23 => "0101010",
		24 => "1111111",
		25 => "1111111",

		26 => "0100001",
		27 => "0100001",	
		28 => "1111111",

		29 => "1111111",
		30 => "1111111",
		31 => "1111111",
		32 => "1111111",

----------part 2---------------

		47 => "1111111",
		48 => "1111110",
		49 => "1111111",

		50 => "0011001",
		51 => "0011001",
		52 => "1111111",
		53 => "1111111",

		54 => "0010001",
		55 => "0011001",
		56 => "1111111",
		57 => "1111111",
	
		58 => "1111111",
		59 => "0001010",
		60 => "1111111",
		61 => "1111111",
	
		62 => "0101001",
		63 => "0101001",
		64 => "1111111",
		65 => "1111111",

		66 => "0100001",
		67 => "0100001",
		68 => "1111111",

		69 => "1111111",
		70 => "1111111",
		71 => "1111111",
		72 => "1111111",

----------part 3---------------

		87 => "1111111",
		88 => "1111110",
		89 => "1111111",

		90 => "0100001",
		91 => "0100001",
		92 => "1111111",
		93 => "1111111",
	
		94 => "1111111",
		95 => "0010010",
		96 => "1111111",	
		97 => "1111111",

		98 => "0101001",
		99 => "0101001",
		100 => "1111111",
	
		101 => "0100001",
		102 => "0100001",
		103 => "1111111",
	
		104 => "0011001",
		105 => "0011001",
		106 => "1111111",

		107 => "1111111",
		108 => "1111111",
		109 => "1111111",
		110 => "1111111",
		111 => "1111111",
		112 => "1111111",

----------part 4---------------

		127 => "1111111",
		128 => "1111110",
		129 => "1111111",

		130 => "1111111",
		131 => "1111111",
		132 => "0010010",
		133 => "1111111",

		134 => "0001001",
		135 => "0001001",
		136 => "1111111",
	
		137 => "0101001",
		138 => "0101001",
		139 => "1111111",
		140 => "0110001",
   	141 => "0110001",
		142 => "1111111",
	
		143 => "1111111",
		144 => "0101010",
		145 => "1111111",
	
		146 => "1111111",
		147 => "1111111",
		148 => "1111111",
		149 => "1111111",
		150 => "1111111",

----------part 5---------------

		167 => "1111111",
		168 => "1111110",
		169 => "1111111",

		170 => "0100001",
		171 => "0100001",
		172 => "1111111",
	
		173 => "0011001",
		174 => "0011001",
		175 => "1111111",
	
		176 => "0010001",
		177 => "0010001",
		178 => "1111111",
		179 => "1111111",
	
		180 => "1111111",
   	181 => "1111111",
		182 => "0001010",
		183 => "1111111",
		184 => "1111111",
	
   	185 => "1111111",
		186 => "1111111",
		187 => "1111111",
		188 => "1111111",
		189 => "1111111",
	others => "0000000"
	);
constant keta5 : matrix := (	
----------------jingle bells------------------------------
--keta5
----------part 1---------------
		7 => "1111111",
		8 => "1111110",
		9 => "1111111",

		10 => "0011001",
		11 => "0011001",
		12 => "1111111",
	
		13 => "1111111",
		14 => "0011001",
		15 => "1111111",
	
		16 => "0011001",
		17 => "0011001",
		18 => "1111111",
	
		19 => "1111111",
		20 => "0011001",
		21 => "1111111",
	
		22 => "0011001",
		23 => "1111111",
		24 => "1111111",
	
		25 => "0011001",
		26 => "0101001",
		27 => "1111111",
	
		28 => "0001001",
		29 => "0010001",
		30 => "0011101",

----------part 2---------------

		47 => "1111111",
		48 => "1111110",
		49 => "1111111",

		50 => "0100001",
		51 => "0100001",
		52 => "1111111",
	
		53 => "0100001",
		54 => "0100001",
		55 => "1111111",
	
		56 => "0100001",
		57 => "0011001",
		58 => "1111111",
	
		59 => "0011001",
		60 => "0011001",
		61 => "0011001",
		62 => "1111111",
	
		63 => "0011001",
		64 => "0010001",
		65 => "1111111",
	
		66 => "0010001",
		67 => "0010001",
		68 => "1111111",
		69 => "0010001",
		70 => "0101001",

----------part 3---------------

		87 => "1111111",
		88 => "1111110",
		89 => "1111111",

		90 => "0011001",
		91 => "0011001",
		92 => "1111111",
	
		93 => "1111111",
		94 => "0011001",
		97 => "1111111",
	
		95 => "0011001",
		96 => "0011001",
		97 => "1111111",
	
		98 => "1111111",
		99 => "0011001",
		100 => "1111111",
	
		101 => "0011001",
		102 => "0101001",
		103 => "1111111",

   	104 => "0001001",
		105 => "0010001",
		106 => "1111111",

		107 => "1111111",
		108 => "0011001",
		109 => "1111111",
   	110 => "1111111",
	
----------part 4---------------

		127 => "1111111",
		128 => "1111110",
		129 => "1111111",

		130 => "0100001",
		131 => "0100001",
		132 => "1111111",
	
		133 => "0100001",
		134 => "0100001",
		135 => "1111111",
	
		136 => "0100001",
		137 => "0100001",
		138 => "1111111",
	
		139 => "0011001",
		140 => "0011001",
   	141 => "0110001",
	
		142 => "1111111",
		143 => "0101001",
		144 => "0101001",
	
		145 => "1111111",
		146 => "0100001",
		147 => "0010001",
	
		148 => "1111111",	149 => "0001010",	150 => "1111111",
	others => "0000000"
	);

constant keta6 : matrix := (
-------little spider-----------
--keta6
----------part 1---------------

   	7 => "1111111",
		8 => "1111110",
		9 => "1111111",

		10 => "1111111",
		11 => "0101001",
		12 => "1111111",
	
		13 => "0001001",
		14 => "0001001",
		15 => "0001001",
	
		16 => "1111111",
		17 => "0010001",
		18 => "0011001",
	
		19 => "1111111",
		20 => "0011001",
		21 => "1111111",
	
		22 => "1111111",
		23 => "0011001",
		24 => "0010001",
	
		25 => "1111111",
		26 => "0001001",
		27 => "1111111",
		28 => "1111111",
	
		29 => "1111111",
		30 => "0010001",
		31 => "0011001",
		32 => "1111111",
	
		33 => "1111111",
		34 => "1111111",
		35 => "0001001",
		36 => "1111111",
		37 => "1111111",

----------part 2---------------
   	47 => "1111111",
		48 => "1111110",
		49 => "1111111",

		50 => "0011001",
		51 => "0011001",
		52 => "1111111",
	
		53 => "1111111",
		54 => "0100001",
		55 => "1111111",
	
		56 => "0101001",
		57 => "0101001",
		58 => "1111111",
	
		59 => "1111111",
		60 => "0100001",
		61 => "0011001",
		62 => "0100001",
		63 => "0101001",
		64 => "0011001",
		65 => "1111111",

		66 => "0001001",
		67 => "0010001",
		68 => "0010001",

		69 => "0011001",
		70 => "0011001",

----------part 3---------------
   	87 => "1111111",
		88 => "1111110",
		89 => "1111111",

		90 => "0010001",
		91 => "0001001",
		92 => "1111111",
	
		93 => "0010001",
		94 => "0011001",
		95 => "1111111",
	
		96 => "1111111",
		97 => "0011001",
		98 => "1111111",
	
		99 => "0010001",
		100 => "0010001",
		101 => "1111111",
	
		102 => "1111111",
		103 => "0001001",
		104 => "0001001",

   	105 => "1111111",
		106 => "0001001",
		107 => "0010001",

		108 => "1111111",
		109 => "0010001",
		110 => "0011001",

		111 => "1111111",
		112 => "0011001",
		113 => "0011001",
	
		114 => "1111111",
		115 => "1111111",
		116 => "1111111",
		117 => "1111111",

----------part 4---------------

		127 => "1111111",
		128 => "1111110",
		129 => "1111111",

		130 => "1111111",
		131 => "0010001",
		132 => "1111111",
		133 => "1111111",

		134 => "0001001",
		135 => "0010001",
		136 => "1111111",
	
		137 => "1111111",
		138 => "0011001",
	139 => "0001001",
	140 => "1111111",
	others => "0000000"
	);
constant keta7 : matrix := (
---------Bus on the wheels-------
--keta7
----------part 1---------------

   	7 => "1111111" ,
		8 => "1111110" ,
		9 => "1111111" ,

		10 => "1111111" ,
		11 => "0001001" ,
		12 => "1111111" ,
	
		13 => "1111111" ,
		14 => "0100001" ,
		15 => "0100001" ,
	
		16 => "1111111" ,
		17 => "0100001" ,
		18 => "0100001" ,
	
		19 => "1111111" ,
		20 => "0110001" ,
		21 => "1111111" ,
	
		22 => "1111111" ,
		23 => "0111001" ,
		24 => "1111111" ,
	
		25 => "1111111" ,
		26 => "0110001" ,
		27 => "1111111" ,
	
		28 => "1111111" ,
		29 => "0100001" ,
		30 => "1111111" ,

----------part 2---------------

		47 => "1111111" ,
		48 => "1111110" ,
		49 => "1111111" ,
	
		50 => "1111111" ,
		51 => "0101001" ,
		52 => "1111111" ,
	
		53 => "1111111" ,
		54 => "0011001" ,
		55 => "1111111" ,
	
		56 => "1111111" ,
		57 => "0001001" ,	
		58 => "1111111" ,
	
		59 => "1111111" ,
		60 => "1101001" ,
		61 => "1111111" ,
	
		62 => "1111111" ,
		63 => "0110001" ,
		64 => "1111111" ,
	
		65 => "1111111" ,
		66 => "0100001" ,
		67 => "1111111" ,
	
		68 => "1111111" ,
		69 => "1111111" ,
		70 => "1111111" ,



----------part 3---------------
   	87 => "1111111" ,	88 => "1111110" ,	89 => "1111111" ,

		90 => "1111111" ,
		91 => "0001001" ,
		92 => "1111111" ,
	
		93 => "1111111" ,
		94 => "0100001" ,
		95 => "0100001" ,
	
		96 => "1111111" ,
		97 => "0100001" ,
		98 => "0100001" ,
	
		99 => "1111111" ,
		100 => "0110001" ,
		101 => "1111111" ,
	
		102 => "1111111" ,
		103 => "0111001" ,
		104 => "1111111" ,
	
		105 => "1111111" ,
		106 => "0110001" ,
		107 => "1111111" ,
	
		108 => "1111111" ,
		109 => "0100001" ,
		110 => "1111111" ,

----------part 4---------------

		127 => "1111111" ,
		128 => "1111110" ,
		129 => "1111111" ,

		130 => "1111111" ,
		131 => "1111111" ,
		132 => "0101001" ,
		133 => "1111111" ,

		134 => "1111111" ,
		135 => "0001001" ,
		136 => "1111111" ,
	
		137 => "1111111" ,
		138 => "0100001" ,
		139 => "1111111" ,
	others => "0000000"
	);
end package;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity MI1 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_MI1 of MI1 is
begin
	y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000111111111111111111111111111111110000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000011111111111111111111111111111111000000000011000000000000001100000000000000110000000000000011000000000000001100000000001111110000000001111111000000001111111100001111111111111111111111111111111100001111111100000000011111100000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		

end architecture; 


--
--
--
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--1111111111111111
--1111111111111111
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000000000110000
--0000001111110000
--0000011111110000
--0000111111110000
--1111111111111111
--1111111111111111
--0000111111110000
--0000011111100000
--0000001111000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000



library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity lines is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_lines of lines is
begin
	y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		

end architecture; 








--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--1111111111111111
--1111111111111111
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000
--0000000000000000


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity re4 is
port (y:out std_logic_vector(0 to 1023));

end entity;

architecture arch_re4 of re4 is
begin
	y<="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000111100000000000011110000111111111111111111111111111111110000000011001110000000001100111000000000110000100000000011000010000000001111000000000000111100000000000011111100000000001111110011111111111111111111111111111111000000001100001000000000110000100000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000001111111111111111111111111111111100011111110000000011111111000000001111111100000000111111110000000011111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

end architecture; 